`include "alarma_desc_conductual.v"

module Newmodule;
    
    alarma_desc_conductual alarma_desc_conductual(/*AUTOINST*/);
endmodule


