`include "alarma_desc_conductual.v"

module autoinst;
    
<<<<<<< HEAD
    alarma_desc_conductual alarma_desc_conductual(/*AUTOINST*/
						  // Outputs
						  .sAlr			(sAlr),
						  // Inputs
						  .sLuz			(sLuz),
						  .sPrta		(sPrta),
						  .sIgn			(sIgn));
endmodule
=======
    alarma_desc_conductual alarma_desc_conductual(/*AUTOINST*/
						  // Outputs
						  .sAlr			(sAlr),
						  // Inputs
						  .sLuz			(sLuz),
						  .sPrta		(sPrta),
						  .sIgn			(sIgn));
>>>>>>> 9265db3b7bc6f32df36467bbe1d86ad8fa17fc0c

endmodule

